** sch_path: /home/ic_design_trg/lna_ihp/xschem/inv.sch
.subckt inv vdd inp out vss
*.PININFO vss:B out:B inp:B vdd:B
M1 out inp vss vss sg13_lv_nmos w=1.0u l=0.72u ng=1 m=1
M2 out inp vdd vdd sg13_lv_pmos w=1.0u l=0.72u ng=1 m=1
.ends
