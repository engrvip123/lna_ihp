** sch_path: /home/ic_design_trg/lna_ihp/xschem/test_dcsweep.sch
**.subckt test_dcsweep
Vgs G GND 'vg'
Vds D GND 0.5
Vd D net1 0
.save i(vd)
XM1 net1 G GND GND sg13_lv_nmos w=5u l=0.25u ng=1 m=40
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt




.include ~/lna_ihp/xschem/simulations/test_dcsweep.save
.param temp=27 wid=70.0u vg=0.45


.control
save all
save @n.xm1.nsg13_lv_nmos[vds]
save @n.xm1.nsg13_lv_nmos[gds]
save @n.xm1.nsg13_lv_nmos[cgs]
save @n.xm1.nsg13_lv_nmos[cgd]
save @n.xm1.nsg13_lv_nmos[vdsat]


op
write test_dcsweep.raw
set appendwrite

* --- wid = 1u ---
*alterparam wid=1u
alterparam vg=0.4
reset
op
set appendwrite
dc Vds 0 1.2 0.01
write test_dcsweep.raw
set appendwrite


* --- wid = 10u ---
*alterparam wid=10u
alterparam vg=0.5
reset
dc Vds 0 1.2 0.01
write test_dcsweep.raw
set appendwrite


* --- wid = 20u ---
*alterparam wid=20u
alterparam vg=0.6
reset
dc Vds 0 1.2 0.01
write test_dcsweep.raw

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
