* Qucs 25.2.0  /home/ic_design_trg/lna_ihp/qucs/lna_prj/lna.sch
.INCLUDE "/usr/local/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_nmos  gnd d g s b w=0.15u l=0.15u ng=1 m=1 mismatch=0 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.34e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 mlist=1
X1 d g s b  sg13_lv_nmos w={w} l={l} ng={ng} m={m} mm_ok={mismatch} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout} 
.ENDS
  
.SUBCKT ind_lumped _net0 _net1 
L1 _net0 _net2  {LSERIES} 
R1 _net2 _net1  {RSERIES} tc1=0.0 tc2=0.0 
C1 _net3 _net0  {CSHUNT1} 
R2 0 _net3  {RSHUNT1} tc1=0.0 tc2=0.0 
C2 _net4 _net1  {CSHUNT2} 
R3 0 _net4  {RSHUNT2} tc1=0.0 tc2=0.0 
.ENDS
.LIB cornerMOSlv.lib mos_tt

.save all @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[gm]
.save all @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[gds]
.save all @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[cgs]
.save all @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[cgd]
.save all @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[cdb]
.save all @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[vth]
.save all @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[vgs]
.save all @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[ids]

.PARAM Lseries = 10n
.PARAM Rseries = 1
.PARAM Cshunt1 = 100f
.PARAM Rshunt1 = 1k
.PARAM Cshunt2 = 100f
.PARAM Rshunt2 = 1k
V1 vdd  0 1.2
VP1 _net0 0 dc 0 ac 0.632456 SIN(0 0.632456 1MEG) portnum 1 z0 50
R1 _net1 n4  10K tc1=0.0 tc2=0.0 
VP2 _net2 0 dc 0 ac 0.632456 SIN(0 0.632456 1MEG) portnum 2 z0 50
LQ1 vdd _net_LQ1 L='5N'
RLQ1 _net_LQ1 n1 R='8*atan(1)*(5N)*(1100MEG)/(10)'
C2 _net0 n4  20P 

Xsg13_lv_nmos1 0 _net3 n3 n2 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=300U l=0.18U ng=1 m=1 mismatch=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.34E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
LQ2 n4 _net_LQ2 L='20N'
RLQ2 _net_LQ2 n3 R='8*atan(1)*(20N)*(1100MEG)/(10)'
Xsg13_lv_nmos2 0 n1 vdd _net3 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=300U l=0.18U ng=1 m=1 mismatch=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.34E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
V2 _net1 0 DC 0.6
C1 n1 _net2  5P 
XSUB 0 n2 ind_lumped

.control

op
let mos_gm = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[gm]
let mos_gds = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[gds]
let mos_cgs = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[cgs]
let mos_cgd = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[cgd]
let mos_cdb = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[cdb]
let mos_vth = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[vth]
let mos_vgs = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[vgs]
let mos_ids = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[ids]
print v(n1) v(n2) v(n3) v(n4) v(vdd)  mos_gm mos_gds mos_cgs mos_cgd mos_cdb mos_vth mos_vgs mos_ids > spice4qucs.dc1.ngspice.dc.print
destroy all
reset

SP DEC 50 1MEG 5G 1
let db_s11 = dB(S_1_1)
let db_s21 = dB(S_2_1)
let db_s12 = dB(S_1_2)
let db_s22 = dB(S_2_2)
let mos_gm = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[gm]
let mos_gds = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[gds]
let mos_cgs = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[cgs]
let mos_cgd = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[cgd]
let mos_cdb = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[cdb]
let mos_vth = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[vth]
let mos_vgs = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[vgs]
let mos_ids = @n.Xsg13_lv_nmos1.x1.nsg13_lv_nmos[ids]
write spice4qucs.sp1.plot S_1_1 Y_1_1 Z_1_1 Cy_1_1 S_1_2 Y_1_2 Z_1_2 Cy_1_2 S_2_1 Y_2_1 Z_2_1 Cy_2_1 S_2_2 Y_2_2 Z_2_2 Cy_2_2 Rn NF SOpt NFmin db_s11 db_s21 db_s12 db_s22 mos_gm mos_gds mos_cgs mos_cgd mos_cdb mos_vth mos_vgs mos_ids
destroy all
reset

exit
.endc
.END
