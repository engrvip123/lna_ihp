** sch_path: /home/ic_design_trg/lna_ihp/xschem/inv_tb.sch
**.subckt inv_tb
Vin in GND dc 0 ac 0 pulse(0, 1.2, 0, 100p, 100p, 2n, 4n )
Vdd net1 GND 1.2
x1 net1 in out GND inv
C1 out GND 1p m=1
**** begin user architecture code


.param temp=27
.control
save all
tran 0.1n 100n
meas tran tdelay TRIG v(in) VAl=0.9 FALl=1 TARG v(out) VAl=0.9 RISE=1
write inv.raw
.endc



.lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/ic_design_trg/lna_ihp/xschem/inv.sym
** sch_path: /home/ic_design_trg/lna_ihp/xschem/inv.sch
.subckt inv vdd inp out vss
*.iopin vss
*.iopin out
*.iopin inp
*.iopin vdd
XM1 out inp vss vss sg13_lv_nmos w=1.0u l=0.72u ng=1 m=1 rfmode=1
XM2 out inp vdd vdd sg13_lv_pmos w=5.0u l=0.72u ng=1 m=1 rfmode=1
.ends

.GLOBAL GND
.end
