** sch_path: /home/ic_design_trg/lna_ihp/xschem/phs_nmos.sch
**.subckt phs_nmos rf_out
*.iopin rf_out
V2 b0 GND b0
V3 b1 GND b1
V4 b2 GND b2
V5 b3 GND b3
V6 b4 GND b4
L8 rf_inp rf_out 6n m=1
C6 rf_out n0 0.2p m=1
C7 rf_out n1 0.4p m=1
C8 rf_out n2 0.8p m=1
C9 rf_out n3 1.6p m=1
C10 rf_out n4 3.2p m=1
V7 rf_inp GND DC 0 AC 1
XM5 n0 b0 GND GND sg13_lv_nmos w=10u l=0.13u ng=1 m=10
XM7 n1 b1 GND GND sg13_lv_nmos w=10u l=0.13u ng=1 m=10
XM8 n2 b2 GND GND sg13_lv_nmos w=10u l=0.13u ng=1 m=10
XM9 n3 b3 GND GND sg13_lv_nmos w=10u l=0.13u ng=1 m=10
XM10 n4 b4 GND GND sg13_lv_nmos w=10u l=0.13u ng=1 m=10
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.param temp=27
.control
save all
save vp(rf_out)

op
write phs_nmos.raw
setappendwrite

ac dec 101 10e6 10e9
meas ac ph_rfout FIND vp(rf_out) AT=1.1182G
meas ac mag_rfout FIND vm(rf_out) AT=1.1182G
write phs_nmos.raw

.endc





.param
+ b0=1.2
+ b1=0
+ b2=0
+ b3=0
+ b4=0


**** end user architecture code
**.ends
.GLOBAL GND
.end
