** sch_path: /home/ic_design_trg/pdk/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/ac_mim_cap.sch
**.subckt ac_mim_cap
V1 in GND dc 0 ac 1
R2 out GND 100k m=1
XC1 out in cap_cmim w=10.0e-6 l=70.0e-6 m=1
**** begin user architecture code



.control
save all
ac dec 1000 1e6 1e9
let mag=abs(out)
meas ac freq_at when mag = 0.707
let C = 1/(2*PI*freq_at*1e+5)
print C
write ac_mim_cap.raw
.endc



.lib /home/ic_design_trg/pdk/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ

**** end user architecture code
**.ends
.GLOBAL GND
.end
