.subckt inv VDD VSS
.ends
.end
